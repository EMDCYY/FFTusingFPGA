library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity TestData is
port(
     clk : in  std_logic;
	  num : in  Std_logic_vector(9 DOWNTO 0) := "0000000000";
	  da1 : out std_logic_vector(11 downto 0);
     da2 : out std_logic_vector(11 downto 0)	  
	  );
end TestData;

architecture Behavioral of TestData is
signal number : integer range 0 to 1024;

TYPE matrix_index is array (0 to 1023) of std_logic_vector(11 downto 0);
--constant R1 : matrix_index :=(
--"100000000000",
--"100000010010",
--"100000100100",
--"100000110110",
--"100001001000",
--"100001011010",
--"100001101100",
--"100001111110",
--"100010001111",
--"100010100001",
--"100010110011",
--"100011000100",
--"100011010110",
--"100011100111",
--"100011111000",
--"100100001001",
--"100100011010",
--"100100101010",
--"100100111011",
--"100101001011",
--"100101011011",
--"100101101011",
--"100101111011",
--"100110001010",
--"100110011001",
--"100110101000",
--"100110110111",
--"100111000101",
--"100111010011",
--"100111100001",
--"100111101111",
--"100111111100",
--"101000001001",
--"101000010101",
--"101000100010",
--"101000101110",
--"101000111001",
--"101001000101",
--"101001010000",
--"101001011010",
--"101001100101",
--"101001101110",
--"101001111000",
--"101010000001",
--"101010001010",
--"101010010010",
--"101010011010",
--"101010100010",
--"101010101001",
--"101010101111",
--"101010110110",
--"101010111100",
--"101011000001",
--"101011000110",
--"101011001011",
--"101011001111",
--"101011010011",
--"101011010110",
--"101011011001",
--"101011011011",
--"101011011101",
--"101011011111",
--"101011100000",
--"101011100001",
--"101011100001",
--"101011100001",
--"101011100000",
--"101011011111",
--"101011011101",
--"101011011011",
--"101011011001",
--"101011010110",
--"101011010011",
--"101011001111",
--"101011001011",
--"101011000110",
--"101011000001",
--"101010111100",
--"101010110110",
--"101010101111",
--"101010101001",
--"101010100010",
--"101010011010",
--"101010010010",
--"101010001010",
--"101010000001",
--"101001111000",
--"101001101110",
--"101001100101",
--"101001011010",
--"101001010000",
--"101001000101",
--"101000111001",
--"101000101110",
--"101000100010",
--"101000010101",
--"101000001001",
--"100111111100",
--"100111101111",
--"100111100001",
--"100111010011",
--"100111000101",
--"100110110111",
--"100110101000",
--"100110011001",
--"100110001010",
--"100101111011",
--"100101101011",
--"100101011011",
--"100101001011",
--"100100111011",
--"100100101010",
--"100100011010",
--"100100001001",
--"100011111000",
--"100011100111",
--"100011010110",
--"100011000100",
--"100010110011",
--"100010100001",
--"100010001111",
--"100001111110",
--"100001101100",
--"100001011010",
--"100001001000",
--"100000110110",
--"100000100100",
--"100000010010",
--"100000000000",
--"011111101101",
--"011111011011",
--"011111001001",
--"011110110111",
--"011110100101",
--"011110010011",
--"011110000001",
--"011101110000",
--"011101011110",
--"011101001100",
--"011100111011",
--"011100101001",
--"011100011000",
--"011100000111",
--"011011110110",
--"011011100101",
--"011011010101",
--"011011000100",
--"011010110100",
--"011010100100",
--"011010010100",
--"011010000100",
--"011001110101",
--"011001100110",
--"011001010111",
--"011001001000",
--"011000111010",
--"011000101100",
--"011000011110",
--"011000010000",
--"011000000011",
--"010111110110",
--"010111101010",
--"010111011101",
--"010111010001",
--"010111000110",
--"010110111010",
--"010110101111",
--"010110100101",
--"010110011010",
--"010110010001",
--"010110000111",
--"010101111110",
--"010101110101",
--"010101101101",
--"010101100101",
--"010101011101",
--"010101010110",
--"010101010000",
--"010101001001",
--"010101000011",
--"010100111110",
--"010100111001",
--"010100110100",
--"010100110000",
--"010100101100",
--"010100101001",
--"010100100110",
--"010100100100",
--"010100100010",
--"010100100000",
--"010100011111",
--"010100011110",
--"010100011110",
--"010100011110",
--"010100011111",
--"010100100000",
--"010100100010",
--"010100100100",
--"010100100110",
--"010100101001",
--"010100101100",
--"010100110000",
--"010100110100",
--"010100111001",
--"010100111110",
--"010101000011",
--"010101001001",
--"010101010000",
--"010101010110",
--"010101011101",
--"010101100101",
--"010101101101",
--"010101110101",
--"010101111110",
--"010110000111",
--"010110010001",
--"010110011010",
--"010110100101",
--"010110101111",
--"010110111010",
--"010111000110",
--"010111010001",
--"010111011101",
--"010111101010",
--"010111110110",
--"011000000011",
--"011000010000",
--"011000011110",
--"011000101100",
--"011000111010",
--"011001001000",
--"011001010111",
--"011001100110",
--"011001110101",
--"011010000100",
--"011010010100",
--"011010100100",
--"011010110100",
--"011011000100",
--"011011010101",
--"011011100101",
--"011011110110",
--"011100000111",
--"011100011000",
--"011100101001",
--"011100111011",
--"011101001100",
--"011101011110",
--"011101110000",
--"011110000001",
--"011110010011",
--"011110100101",
--"011110110111",
--"011111001001",
--"011111011011",
--"011111101101",
--"100000000000",
--"100000010010",
--"100000100100",
--"100000110110",
--"100001001000",
--"100001011010",
--"100001101100",
--"100001111110",
--"100010001111",
--"100010100001",
--"100010110011",
--"100011000100",
--"100011010110",
--"100011100111",
--"100011111000",
--"100100001001",
--"100100011010",
--"100100101010",
--"100100111011",
--"100101001011",
--"100101011011",
--"100101101011",
--"100101111011",
--"100110001010",
--"100110011001",
--"100110101000",
--"100110110111",
--"100111000101",
--"100111010011",
--"100111100001",
--"100111101111",
--"100111111100",
--"101000001001",
--"101000010101",
--"101000100010",
--"101000101110",
--"101000111001",
--"101001000101",
--"101001010000",
--"101001011010",
--"101001100101",
--"101001101110",
--"101001111000",
--"101010000001",
--"101010001010",
--"101010010010",
--"101010011010",
--"101010100010",
--"101010101001",
--"101010101111",
--"101010110110",
--"101010111100",
--"101011000001",
--"101011000110",
--"101011001011",
--"101011001111",
--"101011010011",
--"101011010110",
--"101011011001",
--"101011011011",
--"101011011101",
--"101011011111",
--"101011100000",
--"101011100001",
--"101011100001",
--"101011100001",
--"101011100000",
--"101011011111",
--"101011011101",
--"101011011011",
--"101011011001",
--"101011010110",
--"101011010011",
--"101011001111",
--"101011001011",
--"101011000110",
--"101011000001",
--"101010111100",
--"101010110110",
--"101010101111",
--"101010101001",
--"101010100010",
--"101010011010",
--"101010010010",
--"101010001010",
--"101010000001",
--"101001111000",
--"101001101110",
--"101001100101",
--"101001011010",
--"101001010000",
--"101001000101",
--"101000111001",
--"101000101110",
--"101000100010",
--"101000010101",
--"101000001001",
--"100111111100",
--"100111101111",
--"100111100001",
--"100111010011",
--"100111000101",
--"100110110111",
--"100110101000",
--"100110011001",
--"100110001010",
--"100101111011",
--"100101101011",
--"100101011011",
--"100101001011",
--"100100111011",
--"100100101010",
--"100100011010",
--"100100001001",
--"100011111000",
--"100011100111",
--"100011010110",
--"100011000100",
--"100010110011",
--"100010100001",
--"100010001111",
--"100001111110",
--"100001101100",
--"100001011010",
--"100001001000",
--"100000110110",
--"100000100100",
--"100000010010",
--"100000000000",
--"011111101101",
--"011111011011",
--"011111001001",
--"011110110111",
--"011110100101",
--"011110010011",
--"011110000001",
--"011101110000",
--"011101011110",
--"011101001100",
--"011100111011",
--"011100101001",
--"011100011000",
--"011100000111",
--"011011110110",
--"011011100101",
--"011011010101",
--"011011000100",
--"011010110100",
--"011010100100",
--"011010010100",
--"011010000100",
--"011001110101",
--"011001100110",
--"011001010111",
--"011001001000",
--"011000111010",
--"011000101100",
--"011000011110",
--"011000010000",
--"011000000011",
--"010111110110",
--"010111101010",
--"010111011101",
--"010111010001",
--"010111000110",
--"010110111010",
--"010110101111",
--"010110100101",
--"010110011010",
--"010110010001",
--"010110000111",
--"010101111110",
--"010101110101",
--"010101101101",
--"010101100101",
--"010101011101",
--"010101010110",
--"010101010000",
--"010101001001",
--"010101000011",
--"010100111110",
--"010100111001",
--"010100110100",
--"010100110000",
--"010100101100",
--"010100101001",
--"010100100110",
--"010100100100",
--"010100100010",
--"010100100000",
--"010100011111",
--"010100011110",
--"010100011110",
--"010100011110",
--"010100011111",
--"010100100000",
--"010100100010",
--"010100100100",
--"010100100110",
--"010100101001",
--"010100101100",
--"010100110000",
--"010100110100",
--"010100111001",
--"010100111110",
--"010101000011",
--"010101001001",
--"010101010000",
--"010101010110",
--"010101011101",
--"010101100101",
--"010101101101",
--"010101110101",
--"010101111110",
--"010110000111",
--"010110010001",
--"010110011010",
--"010110100101",
--"010110101111",
--"010110111010",
--"010111000110",
--"010111010001",
--"010111011101",
--"010111101010",
--"010111110110",
--"011000000011",
--"011000010000",
--"011000011110",
--"011000101100",
--"011000111010",
--"011001001000",
--"011001010111",
--"011001100110",
--"011001110101",
--"011010000100",
--"011010010100",
--"011010100100",
--"011010110100",
--"011011000100",
--"011011010101",
--"011011100101",
--"011011110110",
--"011100000111",
--"011100011000",
--"011100101001",
--"011100111011",
--"011101001100",
--"011101011110",
--"011101110000",
--"011110000001",
--"011110010011",
--"011110100101",
--"011110110111",
--"011111001001",
--"011111011011",
--"011111101101",
--"011111111111",
--"100000010010",
--"100000100100",
--"100000110110",
--"100001001000",
--"100001011010",
--"100001101100",
--"100001111110",
--"100010001111",
--"100010100001",
--"100010110011",
--"100011000100",
--"100011010110",
--"100011100111",
--"100011111000",
--"100100001001",
--"100100011010",
--"100100101010",
--"100100111011",
--"100101001011",
--"100101011011",
--"100101101011",
--"100101111011",
--"100110001010",
--"100110011001",
--"100110101000",
--"100110110111",
--"100111000101",
--"100111010011",
--"100111100001",
--"100111101111",
--"100111111100",
--"101000001001",
--"101000010101",
--"101000100010",
--"101000101110",
--"101000111001",
--"101001000101",
--"101001010000",
--"101001011010",
--"101001100101",
--"101001101110",
--"101001111000",
--"101010000001",
--"101010001010",
--"101010010010",
--"101010011010",
--"101010100010",
--"101010101001",
--"101010101111",
--"101010110110",
--"101010111100",
--"101011000001",
--"101011000110",
--"101011001011",
--"101011001111",
--"101011010011",
--"101011010110",
--"101011011001",
--"101011011011",
--"101011011101",
--"101011011111",
--"101011100000",
--"101011100001",
--"101011100001",
--"101011100001",
--"101011100000",
--"101011011111",
--"101011011101",
--"101011011011",
--"101011011001",
--"101011010110",
--"101011010011",
--"101011001111",
--"101011001011",
--"101011000110",
--"101011000001",
--"101010111100",
--"101010110110",
--"101010101111",
--"101010101001",
--"101010100010",
--"101010011010",
--"101010010010",
--"101010001010",
--"101010000001",
--"101001111000",
--"101001101110",
--"101001100101",
--"101001011010",
--"101001010000",
--"101001000101",
--"101000111001",
--"101000101110",
--"101000100010",
--"101000010101",
--"101000001001",
--"100111111100",
--"100111101111",
--"100111100001",
--"100111010011",
--"100111000101",
--"100110110111",
--"100110101000",
--"100110011001",
--"100110001010",
--"100101111011",
--"100101101011",
--"100101011011",
--"100101001011",
--"100100111011",
--"100100101010",
--"100100011010",
--"100100001001",
--"100011111000",
--"100011100111",
--"100011010110",
--"100011000100",
--"100010110011",
--"100010100001",
--"100010001111",
--"100001111110",
--"100001101100",
--"100001011010",
--"100001001000",
--"100000110110",
--"100000100100",
--"100000010010",
--"100000000000",
--"011111101101",
--"011111011011",
--"011111001001",
--"011110110111",
--"011110100101",
--"011110010011",
--"011110000001",
--"011101110000",
--"011101011110",
--"011101001100",
--"011100111011",
--"011100101001",
--"011100011000",
--"011100000111",
--"011011110110",
--"011011100101",
--"011011010101",
--"011011000100",
--"011010110100",
--"011010100100",
--"011010010100",
--"011010000100",
--"011001110101",
--"011001100110",
--"011001010111",
--"011001001000",
--"011000111010",
--"011000101100",
--"011000011110",
--"011000010000",
--"011000000011",
--"010111110110",
--"010111101010",
--"010111011101",
--"010111010001",
--"010111000110",
--"010110111010",
--"010110101111",
--"010110100101",
--"010110011010",
--"010110010001",
--"010110000111",
--"010101111110",
--"010101110101",
--"010101101101",
--"010101100101",
--"010101011101",
--"010101010110",
--"010101010000",
--"010101001001",
--"010101000011",
--"010100111110",
--"010100111001",
--"010100110100",
--"010100110000",
--"010100101100",
--"010100101001",
--"010100100110",
--"010100100100",
--"010100100010",
--"010100100000",
--"010100011111",
--"010100011110",
--"010100011110",
--"010100011110",
--"010100011111",
--"010100100000",
--"010100100010",
--"010100100100",
--"010100100110",
--"010100101001",
--"010100101100",
--"010100110000",
--"010100110100",
--"010100111001",
--"010100111110",
--"010101000011",
--"010101001001",
--"010101010000",
--"010101010110",
--"010101011101",
--"010101100101",
--"010101101101",
--"010101110101",
--"010101111110",
--"010110000111",
--"010110010001",
--"010110011010",
--"010110100101",
--"010110101111",
--"010110111010",
--"010111000110",
--"010111010001",
--"010111011101",
--"010111101010",
--"010111110110",
--"011000000011",
--"011000010000",
--"011000011110",
--"011000101100",
--"011000111010",
--"011001001000",
--"011001010111",
--"011001100110",
--"011001110101",
--"011010000100",
--"011010010100",
--"011010100100",
--"011010110100",
--"011011000100",
--"011011010101",
--"011011100101",
--"011011110110",
--"011100000111",
--"011100011000",
--"011100101001",
--"011100111011",
--"011101001100",
--"011101011110",
--"011101110000",
--"011110000001",
--"011110010011",
--"011110100101",
--"011110110111",
--"011111001001",
--"011111011011",
--"011111101101",
--"011111111111",
--"100000010010",
--"100000100100",
--"100000110110",
--"100001001000",
--"100001011010",
--"100001101100",
--"100001111110",
--"100010001111",
--"100010100001",
--"100010110011",
--"100011000100",
--"100011010110",
--"100011100111",
--"100011111000",
--"100100001001",
--"100100011010",
--"100100101010",
--"100100111011",
--"100101001011",
--"100101011011",
--"100101101011",
--"100101111011",
--"100110001010",
--"100110011001",
--"100110101000",
--"100110110111",
--"100111000101",
--"100111010011",
--"100111100001",
--"100111101111",
--"100111111100",
--"101000001001",
--"101000010101",
--"101000100010",
--"101000101110",
--"101000111001",
--"101001000101",
--"101001010000",
--"101001011010",
--"101001100101",
--"101001101110",
--"101001111000",
--"101010000001",
--"101010001010",
--"101010010010",
--"101010011010",
--"101010100010",
--"101010101001",
--"101010101111",
--"101010110110",
--"101010111100",
--"101011000001",
--"101011000110",
--"101011001011",
--"101011001111",
--"101011010011",
--"101011010110",
--"101011011001",
--"101011011011",
--"101011011101",
--"101011011111",
--"101011100000",
--"101011100001",
--"101011100001",
--"101011100001",
--"101011100000",
--"101011011111",
--"101011011101",
--"101011011011",
--"101011011001",
--"101011010110",
--"101011010011",
--"101011001111",
--"101011001011",
--"101011000110",
--"101011000001",
--"101010111100",
--"101010110110",
--"101010101111",
--"101010101001",
--"101010100010",
--"101010011010",
--"101010010010",
--"101010001010",
--"101010000001",
--"101001111000",
--"101001101110",
--"101001100101",
--"101001011010",
--"101001010000",
--"101001000101",
--"101000111001",
--"101000101110",
--"101000100010",
--"101000010101",
--"101000001001",
--"100111111100",
--"100111101111",
--"100111100001",
--"100111010011",
--"100111000101",
--"100110110111",
--"100110101000",
--"100110011001",
--"100110001010",
--"100101111011",
--"100101101011",
--"100101011011",
--"100101001011",
--"100100111011",
--"100100101010",
--"100100011010",
--"100100001001",
--"100011111000",
--"100011100111",
--"100011010110",
--"100011000100",
--"100010110011",
--"100010100001",
--"100010001111",
--"100001111110",
--"100001101100",
--"100001011010",
--"100001001000",
--"100000110110",
--"100000100100",
--"100000010010",
--"100000000000",
--"011111101101",
--"011111011011",
--"011111001001",
--"011110110111",
--"011110100101",
--"011110010011",
--"011110000001",
--"011101110000",
--"011101011110",
--"011101001100",
--"011100111011",
--"011100101001",
--"011100011000",
--"011100000111",
--"011011110110",
--"011011100101",
--"011011010101",
--"011011000100",
--"011010110100",
--"011010100100",
--"011010010100",
--"011010000100",
--"011001110101",
--"011001100110",
--"011001010111",
--"011001001000",
--"011000111010",
--"011000101100",
--"011000011110",
--"011000010000",
--"011000000011",
--"010111110110",
--"010111101010",
--"010111011101",
--"010111010001",
--"010111000110",
--"010110111010",
--"010110101111",
--"010110100101",
--"010110011010",
--"010110010001",
--"010110000111",
--"010101111110",
--"010101110101",
--"010101101101",
--"010101100101",
--"010101011101",
--"010101010110",
--"010101010000",
--"010101001001",
--"010101000011",
--"010100111110",
--"010100111001",
--"010100110100",
--"010100110000",
--"010100101100",
--"010100101001",
--"010100100110",
--"010100100100",
--"010100100010",
--"010100100000",
--"010100011111",
--"010100011110",
--"010100011110",
--"010100011110",
--"010100011111",
--"010100100000",
--"010100100010",
--"010100100100",
--"010100100110",
--"010100101001",
--"010100101100",
--"010100110000",
--"010100110100",
--"010100111001",
--"010100111110",
--"010101000011",
--"010101001001",
--"010101010000",
--"010101010110",
--"010101011101",
--"010101100101",
--"010101101101",
--"010101110101",
--"010101111110",
--"010110000111",
--"010110010001",
--"010110011010",
--"010110100101",
--"010110101111",
--"010110111010",
--"010111000110",
--"010111010001",
--"010111011101",
--"010111101010",
--"010111110110",
--"011000000011",
--"011000010000",
--"011000011110",
--"011000101100",
--"011000111010",
--"011001001000",
--"011001010111",
--"011001100110",
--"011001110101",
--"011010000100",
--"011010010100",
--"011010100100",
--"011010110100",
--"011011000100",
--"011011010101",
--"011011100101",
--"011011110110",
--"011100000111",
--"011100011000",
--"011100101001",
--"011100111011",
--"011101001100",
--"011101011110",
--"011101110000",
--"011110000001",
--"011110010011",
--"011110100101",
--"011110110111",
--"011111001001",
--"011111011011",
--"011111101101"
--);

--constant R2 : matrix_index :=(
--"101000001001",
--"101000010101",
--"101000100010",
--"101000101110",
--"101000111001",
--"101001000101",
--"101001010000",
--"101001011010",
--"101001100101",
--"101001101110",
--"101001111000",
--"101010000001",
--"101010001010",
--"101010010010",
--"101010011010",
--"101010100010",
--"101010101001",
--"101010101111",
--"101010110110",
--"101010111100",
--"101011000001",
--"101011000110",
--"101011001011",
--"101011001111",
--"101011010011",
--"101011010110",
--"101011011001",
--"101011011011",
--"101011011101",
--"101011011111",
--"101011100000",
--"101011100001",
--"101011100001",
--"101011100001",
--"101011100000",
--"101011011111",
--"101011011101",
--"101011011011",
--"101011011001",
--"101011010110",
--"101011010011",
--"101011001111",
--"101011001011",
--"101011000110",
--"101011000001",
--"101010111100",
--"101010110110",
--"101010101111",
--"101010101001",
--"101010100010",
--"101010011010",
--"101010010010",
--"101010001010",
--"101010000001",
--"101001111000",
--"101001101110",
--"101001100101",
--"101001011010",
--"101001010000",
--"101001000101",
--"101000111001",
--"101000101110",
--"101000100010",
--"101000010101",
--"101000001001",
--"100111111100",
--"100111101111",
--"100111100001",
--"100111010011",
--"100111000101",
--"100110110111",
--"100110101000",
--"100110011001",
--"100110001010",
--"100101111011",
--"100101101011",
--"100101011011",
--"100101001011",
--"100100111011",
--"100100101010",
--"100100011010",
--"100100001001",
--"100011111000",
--"100011100111",
--"100011010110",
--"100011000100",
--"100010110011",
--"100010100001",
--"100010001111",
--"100001111110",
--"100001101100",
--"100001011010",
--"100001001000",
--"100000110110",
--"100000100100",
--"100000010010",
--"100000000000",
--"011111101101",
--"011111011011",
--"011111001001",
--"011110110111",
--"011110100101",
--"011110010011",
--"011110000001",
--"011101110000",
--"011101011110",
--"011101001100",
--"011100111011",
--"011100101001",
--"011100011000",
--"011100000111",
--"011011110110",
--"011011100101",
--"011011010101",
--"011011000100",
--"011010110100",
--"011010100100",
--"011010010100",
--"011010000100",
--"011001110101",
--"011001100110",
--"011001010111",
--"011001001000",
--"011000111010",
--"011000101100",
--"011000011110",
--"011000010000",
--"011000000011",
--"010111110110",
--"010111101010",
--"010111011101",
--"010111010001",
--"010111000110",
--"010110111010",
--"010110101111",
--"010110100101",
--"010110011010",
--"010110010001",
--"010110000111",
--"010101111110",
--"010101110101",
--"010101101101",
--"010101100101",
--"010101011101",
--"010101010110",
--"010101010000",
--"010101001001",
--"010101000011",
--"010100111110",
--"010100111001",
--"010100110100",
--"010100110000",
--"010100101100",
--"010100101001",
--"010100100110",
--"010100100100",
--"010100100010",
--"010100100000",
--"010100011111",
--"010100011110",
--"010100011110",
--"010100011110",
--"010100011111",
--"010100100000",
--"010100100010",
--"010100100100",
--"010100100110",
--"010100101001",
--"010100101100",
--"010100110000",
--"010100110100",
--"010100111001",
--"010100111110",
--"010101000011",
--"010101001001",
--"010101010000",
--"010101010110",
--"010101011101",
--"010101100101",
--"010101101101",
--"010101110101",
--"010101111110",
--"010110000111",
--"010110010001",
--"010110011010",
--"010110100101",
--"010110101111",
--"010110111010",
--"010111000110",
--"010111010001",
--"010111011101",
--"010111101010",
--"010111110110",
--"011000000011",
--"011000010000",
--"011000011110",
--"011000101100",
--"011000111010",
--"011001001000",
--"011001010111",
--"011001100110",
--"011001110101",
--"011010000100",
--"011010010100",
--"011010100100",
--"011010110100",
--"011011000100",
--"011011010101",
--"011011100101",
--"011011110110",
--"011100000111",
--"011100011000",
--"011100101001",
--"011100111011",
--"011101001100",
--"011101011110",
--"011101110000",
--"011110000001",
--"011110010011",
--"011110100101",
--"011110110111",
--"011111001001",
--"011111011011",
--"011111101101",
--"100000000000",
--"100000010010",
--"100000100100",
--"100000110110",
--"100001001000",
--"100001011010",
--"100001101100",
--"100001111110",
--"100010001111",
--"100010100001",
--"100010110011",
--"100011000100",
--"100011010110",
--"100011100111",
--"100011111000",
--"100100001001",
--"100100011010",
--"100100101010",
--"100100111011",
--"100101001011",
--"100101011011",
--"100101101011",
--"100101111011",
--"100110001010",
--"100110011001",
--"100110101000",
--"100110110111",
--"100111000101",
--"100111010011",
--"100111100001",
--"100111101111",
--"100111111100",
--"101000001001",
--"101000010101",
--"101000100010",
--"101000101110",
--"101000111001",
--"101001000101",
--"101001010000",
--"101001011010",
--"101001100101",
--"101001101110",
--"101001111000",
--"101010000001",
--"101010001010",
--"101010010010",
--"101010011010",
--"101010100010",
--"101010101001",
--"101010101111",
--"101010110110",
--"101010111100",
--"101011000001",
--"101011000110",
--"101011001011",
--"101011001111",
--"101011010011",
--"101011010110",
--"101011011001",
--"101011011011",
--"101011011101",
--"101011011111",
--"101011100000",
--"101011100001",
--"101011100001",
--"101011100001",
--"101011100000",
--"101011011111",
--"101011011101",
--"101011011011",
--"101011011001",
--"101011010110",
--"101011010011",
--"101011001111",
--"101011001011",
--"101011000110",
--"101011000001",
--"101010111100",
--"101010110110",
--"101010101111",
--"101010101001",
--"101010100010",
--"101010011010",
--"101010010010",
--"101010001010",
--"101010000001",
--"101001111000",
--"101001101110",
--"101001100101",
--"101001011010",
--"101001010000",
--"101001000101",
--"101000111001",
--"101000101110",
--"101000100010",
--"101000010101",
--"101000001001",
--"100111111100",
--"100111101111",
--"100111100001",
--"100111010011",
--"100111000101",
--"100110110111",
--"100110101000",
--"100110011001",
--"100110001010",
--"100101111011",
--"100101101011",
--"100101011011",
--"100101001011",
--"100100111011",
--"100100101010",
--"100100011010",
--"100100001001",
--"100011111000",
--"100011100111",
--"100011010110",
--"100011000100",
--"100010110011",
--"100010100001",
--"100010001111",
--"100001111110",
--"100001101100",
--"100001011010",
--"100001001000",
--"100000110110",
--"100000100100",
--"100000010010",
--"100000000000",
--"011111101101",
--"011111011011",
--"011111001001",
--"011110110111",
--"011110100101",
--"011110010011",
--"011110000001",
--"011101110000",
--"011101011110",
--"011101001100",
--"011100111011",
--"011100101001",
--"011100011000",
--"011100000111",
--"011011110110",
--"011011100101",
--"011011010101",
--"011011000100",
--"011010110100",
--"011010100100",
--"011010010100",
--"011010000100",
--"011001110101",
--"011001100110",
--"011001010111",
--"011001001000",
--"011000111010",
--"011000101100",
--"011000011110",
--"011000010000",
--"011000000011",
--"010111110110",
--"010111101010",
--"010111011101",
--"010111010001",
--"010111000110",
--"010110111010",
--"010110101111",
--"010110100101",
--"010110011010",
--"010110010001",
--"010110000111",
--"010101111110",
--"010101110101",
--"010101101101",
--"010101100101",
--"010101011101",
--"010101010110",
--"010101010000",
--"010101001001",
--"010101000011",
--"010100111110",
--"010100111001",
--"010100110100",
--"010100110000",
--"010100101100",
--"010100101001",
--"010100100110",
--"010100100100",
--"010100100010",
--"010100100000",
--"010100011111",
--"010100011110",
--"010100011110",
--"010100011110",
--"010100011111",
--"010100100000",
--"010100100010",
--"010100100100",
--"010100100110",
--"010100101001",
--"010100101100",
--"010100110000",
--"010100110100",
--"010100111001",
--"010100111110",
--"010101000011",
--"010101001001",
--"010101010000",
--"010101010110",
--"010101011101",
--"010101100101",
--"010101101101",
--"010101110101",
--"010101111110",
--"010110000111",
--"010110010001",
--"010110011010",
--"010110100101",
--"010110101111",
--"010110111010",
--"010111000110",
--"010111010001",
--"010111011101",
--"010111101010",
--"010111110110",
--"011000000011",
--"011000010000",
--"011000011110",
--"011000101100",
--"011000111010",
--"011001001000",
--"011001010111",
--"011001100110",
--"011001110101",
--"011010000100",
--"011010010100",
--"011010100100",
--"011010110100",
--"011011000100",
--"011011010101",
--"011011100101",
--"011011110110",
--"011100000111",
--"011100011000",
--"011100101001",
--"011100111011",
--"011101001100",
--"011101011110",
--"011101110000",
--"011110000001",
--"011110010011",
--"011110100101",
--"011110110111",
--"011111001001",
--"011111011011",
--"011111101101",
--"011111111111",
--"100000010010",
--"100000100100",
--"100000110110",
--"100001001000",
--"100001011010",
--"100001101100",
--"100001111110",
--"100010001111",
--"100010100001",
--"100010110011",
--"100011000100",
--"100011010110",
--"100011100111",
--"100011111000",
--"100100001001",
--"100100011010",
--"100100101010",
--"100100111011",
--"100101001011",
--"100101011011",
--"100101101011",
--"100101111011",
--"100110001010",
--"100110011001",
--"100110101000",
--"100110110111",
--"100111000101",
--"100111010011",
--"100111100001",
--"100111101111",
--"100111111100",
--"101000001001",
--"101000010101",
--"101000100010",
--"101000101110",
--"101000111001",
--"101001000101",
--"101001010000",
--"101001011010",
--"101001100101",
--"101001101110",
--"101001111000",
--"101010000001",
--"101010001010",
--"101010010010",
--"101010011010",
--"101010100010",
--"101010101001",
--"101010101111",
--"101010110110",
--"101010111100",
--"101011000001",
--"101011000110",
--"101011001011",
--"101011001111",
--"101011010011",
--"101011010110",
--"101011011001",
--"101011011011",
--"101011011101",
--"101011011111",
--"101011100000",
--"101011100001",
--"101011100001",
--"101011100001",
--"101011100000",
--"101011011111",
--"101011011101",
--"101011011011",
--"101011011001",
--"101011010110",
--"101011010011",
--"101011001111",
--"101011001011",
--"101011000110",
--"101011000001",
--"101010111100",
--"101010110110",
--"101010101111",
--"101010101001",
--"101010100010",
--"101010011010",
--"101010010010",
--"101010001010",
--"101010000001",
--"101001111000",
--"101001101110",
--"101001100101",
--"101001011010",
--"101001010000",
--"101001000101",
--"101000111001",
--"101000101110",
--"101000100010",
--"101000010101",
--"101000001001",
--"100111111100",
--"100111101111",
--"100111100001",
--"100111010011",
--"100111000101",
--"100110110111",
--"100110101000",
--"100110011001",
--"100110001010",
--"100101111011",
--"100101101011",
--"100101011011",
--"100101001011",
--"100100111011",
--"100100101010",
--"100100011010",
--"100100001001",
--"100011111000",
--"100011100111",
--"100011010110",
--"100011000100",
--"100010110011",
--"100010100001",
--"100010001111",
--"100001111110",
--"100001101100",
--"100001011010",
--"100001001000",
--"100000110110",
--"100000100100",
--"100000010010",
--"100000000000",
--"011111101101",
--"011111011011",
--"011111001001",
--"011110110111",
--"011110100101",
--"011110010011",
--"011110000001",
--"011101110000",
--"011101011110",
--"011101001100",
--"011100111011",
--"011100101001",
--"011100011000",
--"011100000111",
--"011011110110",
--"011011100101",
--"011011010101",
--"011011000100",
--"011010110100",
--"011010100100",
--"011010010100",
--"011010000100",
--"011001110101",
--"011001100110",
--"011001010111",
--"011001001000",
--"011000111010",
--"011000101100",
--"011000011110",
--"011000010000",
--"011000000011",
--"010111110110",
--"010111101010",
--"010111011101",
--"010111010001",
--"010111000110",
--"010110111010",
--"010110101111",
--"010110100101",
--"010110011010",
--"010110010001",
--"010110000111",
--"010101111110",
--"010101110101",
--"010101101101",
--"010101100101",
--"010101011101",
--"010101010110",
--"010101010000",
--"010101001001",
--"010101000011",
--"010100111110",
--"010100111001",
--"010100110100",
--"010100110000",
--"010100101100",
--"010100101001",
--"010100100110",
--"010100100100",
--"010100100010",
--"010100100000",
--"010100011111",
--"010100011110",
--"010100011110",
--"010100011110",
--"010100011111",
--"010100100000",
--"010100100010",
--"010100100100",
--"010100100110",
--"010100101001",
--"010100101100",
--"010100110000",
--"010100110100",
--"010100111001",
--"010100111110",
--"010101000011",
--"010101001001",
--"010101010000",
--"010101010110",
--"010101011101",
--"010101100101",
--"010101101101",
--"010101110101",
--"010101111110",
--"010110000111",
--"010110010001",
--"010110011010",
--"010110100101",
--"010110101111",
--"010110111010",
--"010111000110",
--"010111010001",
--"010111011101",
--"010111101010",
--"010111110110",
--"011000000011",
--"011000010000",
--"011000011110",
--"011000101100",
--"011000111010",
--"011001001000",
--"011001010111",
--"011001100110",
--"011001110101",
--"011010000100",
--"011010010100",
--"011010100100",
--"011010110100",
--"011011000100",
--"011011010101",
--"011011100101",
--"011011110110",
--"011100000111",
--"011100011000",
--"011100101001",
--"011100111011",
--"011101001100",
--"011101011110",
--"011101110000",
--"011110000001",
--"011110010011",
--"011110100101",
--"011110110111",
--"011111001001",
--"011111011011",
--"011111101101",
--"011111111111",
--"100000010010",
--"100000100100",
--"100000110110",
--"100001001000",
--"100001011010",
--"100001101100",
--"100001111110",
--"100010001111",
--"100010100001",
--"100010110011",
--"100011000100",
--"100011010110",
--"100011100111",
--"100011111000",
--"100100001001",
--"100100011010",
--"100100101010",
--"100100111011",
--"100101001011",
--"100101011011",
--"100101101011",
--"100101111011",
--"100110001010",
--"100110011001",
--"100110101000",
--"100110110111",
--"100111000101",
--"100111010011",
--"100111100001",
--"100111101111",
--"100111111100",
--"101000001001",
--"101000010101",
--"101000100010",
--"101000101110",
--"101000111001",
--"101001000101",
--"101001010000",
--"101001011010",
--"101001100101",
--"101001101110",
--"101001111000",
--"101010000001",
--"101010001010",
--"101010010010",
--"101010011010",
--"101010100010",
--"101010101001",
--"101010101111",
--"101010110110",
--"101010111100",
--"101011000001",
--"101011000110",
--"101011001011",
--"101011001111",
--"101011010011",
--"101011010110",
--"101011011001",
--"101011011011",
--"101011011101",
--"101011011111",
--"101011100000",
--"101011100001",
--"101011100001",
--"101011100001",
--"101011100000",
--"101011011111",
--"101011011101",
--"101011011011",
--"101011011001",
--"101011010110",
--"101011010011",
--"101011001111",
--"101011001011",
--"101011000110",
--"101011000001",
--"101010111100",
--"101010110110",
--"101010101111",
--"101010101001",
--"101010100010",
--"101010011010",
--"101010010010",
--"101010001010",
--"101010000001",
--"101001111000",
--"101001101110",
--"101001100101",
--"101001011010",
--"101001010000",
--"101001000101",
--"101000111001",
--"101000101110",
--"101000100010",
--"101000010101",
--"101000001001",
--"100111111100",
--"100111101111",
--"100111100001",
--"100111010011",
--"100111000101",
--"100110110111",
--"100110101000",
--"100110011001",
--"100110001010",
--"100101111011",
--"100101101011",
--"100101011011",
--"100101001011",
--"100100111011",
--"100100101010",
--"100100011010",
--"100100001001",
--"100011111000",
--"100011100111",
--"100011010110",
--"100011000100",
--"100010110011",
--"100010100001",
--"100010001111",
--"100001111110",
--"100001101100",
--"100001011010",
--"100001001000",
--"100000110110",
--"100000100100",
--"100000010010",
--"100000000000",
--"011111101101",
--"011111011011",
--"011111001001",
--"011110110111",
--"011110100101",
--"011110010011",
--"011110000001",
--"011101110000",
--"011101011110",
--"011101001100",
--"011100111011",
--"011100101001",
--"011100011000",
--"011100000111",
--"011011110110",
--"011011100101",
--"011011010101",
--"011011000100",
--"011010110100",
--"011010100100",
--"011010010100",
--"011010000100",
--"011001110101",
--"011001100110",
--"011001010111",
--"011001001000",
--"011000111010",
--"011000101100",
--"011000011110",
--"011000010000",
--"011000000011",
--"010111110110",
--"010111101010",
--"010111011101",
--"010111010001",
--"010111000110",
--"010110111010",
--"010110101111",
--"010110100101",
--"010110011010",
--"010110010001",
--"010110000111",
--"010101111110",
--"010101110101",
--"010101101101",
--"010101100101",
--"010101011101",
--"010101010110",
--"010101010000",
--"010101001001",
--"010101000011",
--"010100111110",
--"010100111001",
--"010100110100",
--"010100110000",
--"010100101100",
--"010100101001",
--"010100100110",
--"010100100100",
--"010100100010",
--"010100100000",
--"010100011111",
--"010100011110",
--"010100011110",
--"010100011110",
--"010100011111",
--"010100100000",
--"010100100010",
--"010100100100",
--"010100100110",
--"010100101001",
--"010100101100",
--"010100110000",
--"010100110100",
--"010100111001",
--"010100111110",
--"010101000011",
--"010101001001",
--"010101010000",
--"010101010110",
--"010101011101",
--"010101100101",
--"010101101101",
--"010101110101",
--"010101111110",
--"010110000111",
--"010110010001",
--"010110011010",
--"010110100101",
--"010110101111",
--"010110111010",
--"010111000110",
--"010111010001",
--"010111011101",
--"010111101010",
--"010111110110",
--"011000000011",
--"011000010000",
--"011000011110",
--"011000101100",
--"011000111010",
--"011001001000",
--"011001010111",
--"011001100110",
--"011001110101",
--"011010000100",
--"011010010100",
--"011010100100",
--"011010110100",
--"011011000100",
--"011011010101",
--"011011100101",
--"011011110110",
--"011100000111",
--"011100011000",
--"011100101001",
--"011100111011",
--"011101001100",
--"011101011110",
--"011101110000",
--"011110000001",
--"011110010011",
--"011110100101",
--"011110110111",
--"011111001001",
--"011111011011",
--"011111101101",
--"100000000000",
--"100000010010",
--"100000100100",
--"100000110110",
--"100001001000",
--"100001011010",
--"100001101100",
--"100001111110",
--"100010001111",
--"100010100001",
--"100010110011",
--"100011000100",
--"100011010110",
--"100011100111",
--"100011111000",
--"100100001001",
--"100100011010",
--"100100101010",
--"100100111011",
--"100101001011",
--"100101011011",
--"100101101011",
--"100101111011",
--"100110001010",
--"100110011001",
--"100110101000",
--"100110110111",
--"100111000101",
--"100111010011",
--"100111100001",
--"100111101111",
--"100111111100"
--);

constant R1 : matrix_index :=(
"110101001011",
"110101101110",
"110110001111",
"110110110000",
"110111010000",
"110111101111",
"111000001101",
"111000101011",
"111001000111",
"111001100010",
"111001111101",
"111010010110",
"111010101110",
"111011000101",
"111011011100",
"111011110001",
"111100000101",
"111100011000",
"111100101010",
"111100111011",
"111101001010",
"111101011001",
"111101100110",
"111101110011",
"111101111110",
"111110001000",
"111110010001",
"111110011000",
"111110011111",
"111110100100",
"111110101000",
"111110101011",
"111110101101",
"111110101110",
"111110101101",
"111110101011",
"111110101000",
"111110100100",
"111110011111",
"111110011000",
"111110010001",
"111110001000",
"111101111110",
"111101110011",
"111101100110",
"111101011001",
"111101001010",
"111100111011",
"111100101010",
"111100011000",
"111100000101",
"111011110001",
"111011011100",
"111011000101",
"111010101110",
"111010010110",
"111001111101",
"111001100010",
"111001000111",
"111000101011",
"111000001101",
"110111101111",
"110111010000",
"110110110000",
"110110001111",
"110101101110",
"110101001011",
"110100101000",
"110100000100",
"110011011111",
"110010111001",
"110010010011",
"110001101100",
"110001000100",
"110000011011",
"101111110010",
"101111001001",
"101110011110",
"101101110011",
"101101001000",
"101100011100",
"101011110000",
"101011000011",
"101010010110",
"101001101000",
"101000111010",
"101000001100",
"100111011101",
"100110101110",
"100101111111",
"100101010000",
"100100100000",
"100011110000",
"100011000000",
"100010010000",
"100001100000",
"100000110000",
"100000000000",
"011111001111",
"011110011111",
"011101101111",
"011100111111",
"011100001111",
"011011011111",
"011010101111",
"011010000000",
"011001010001",
"011000100010",
"010111110011",
"010111000101",
"010110010111",
"010101101001",
"010100111100",
"010100001111",
"010011100011",
"010010110111",
"010010001100",
"010001100001",
"010000110110",
"010000001101",
"001111100100",
"001110111011",
"001110010011",
"001101101100",
"001101000110",
"001100100000",
"001011111011",
"001011010111",
"001010110100",
"001010010001",
"001001110000",
"001001001111",
"001000101111",
"001000010000",
"000111110010",
"000111010100",
"000110111000",
"000110011101",
"000110000010",
"000101101001",
"000101010001",
"000100111010",
"000100100011",
"000100001110",
"000011111010",
"000011100111",
"000011010101",
"000011000100",
"000010110101",
"000010100110",
"000010011001",
"000010001100",
"000010000001",
"000001110111",
"000001101110",
"000001100111",
"000001100000",
"000001011011",
"000001010111",
"000001010100",
"000001010010",
"000001010001",
"000001010010",
"000001010100",
"000001010111",
"000001011011",
"000001100000",
"000001100111",
"000001101110",
"000001110111",
"000010000001",
"000010001100",
"000010011001",
"000010100110",
"000010110101",
"000011000100",
"000011010101",
"000011100111",
"000011111010",
"000100001110",
"000100100011",
"000100111010",
"000101010001",
"000101101001",
"000110000010",
"000110011101",
"000110111000",
"000111010100",
"000111110010",
"001000010000",
"001000101111",
"001001001111",
"001001110000",
"001010010001",
"001010110100",
"001011010111",
"001011111011",
"001100100000",
"001101000110",
"001101101100",
"001110010011",
"001110111011",
"001111100100",
"010000001101",
"010000110110",
"010001100001",
"010010001100",
"010010110111",
"010011100011",
"010100001111",
"010100111100",
"010101101001",
"010110010111",
"010111000101",
"010111110011",
"011000100010",
"011001010001",
"011010000000",
"011010101111",
"011011011111",
"011100001111",
"011100111111",
"011101101111",
"011110011111",
"011111001111",
"011111111111",
"100000110000",
"100001100000",
"100010010000",
"100011000000",
"100011110000",
"100100100000",
"100101010000",
"100101111111",
"100110101110",
"100111011101",
"101000001100",
"101000111010",
"101001101000",
"101010010110",
"101011000011",
"101011110000",
"101100011100",
"101101001000",
"101101110011",
"101110011110",
"101111001001",
"101111110010",
"110000011011",
"110001000100",
"110001101100",
"110010010011",
"110010111001",
"110011011111",
"110100000100",
"110100101000",
"110101001011",
"110101101110",
"110110001111",
"110110110000",
"110111010000",
"110111101111",
"111000001101",
"111000101011",
"111001000111",
"111001100010",
"111001111101",
"111010010110",
"111010101110",
"111011000101",
"111011011100",
"111011110001",
"111100000101",
"111100011000",
"111100101010",
"111100111011",
"111101001010",
"111101011001",
"111101100110",
"111101110011",
"111101111110",
"111110001000",
"111110010001",
"111110011000",
"111110011111",
"111110100100",
"111110101000",
"111110101011",
"111110101101",
"111110101110",
"111110101101",
"111110101011",
"111110101000",
"111110100100",
"111110011111",
"111110011000",
"111110010001",
"111110001000",
"111101111110",
"111101110011",
"111101100110",
"111101011001",
"111101001010",
"111100111011",
"111100101010",
"111100011000",
"111100000101",
"111011110001",
"111011011100",
"111011000101",
"111010101110",
"111010010110",
"111001111101",
"111001100010",
"111001000111",
"111000101011",
"111000001101",
"110111101111",
"110111010000",
"110110110000",
"110110001111",
"110101101110",
"110101001011",
"110100101000",
"110100000100",
"110011011111",
"110010111001",
"110010010011",
"110001101100",
"110001000100",
"110000011011",
"101111110010",
"101111001001",
"101110011110",
"101101110011",
"101101001000",
"101100011100",
"101011110000",
"101011000011",
"101010010110",
"101001101000",
"101000111010",
"101000001100",
"100111011101",
"100110101110",
"100101111111",
"100101010000",
"100100100000",
"100011110000",
"100011000000",
"100010010000",
"100001100000",
"100000110000",
"100000000000",
"011111001111",
"011110011111",
"011101101111",
"011100111111",
"011100001111",
"011011011111",
"011010101111",
"011010000000",
"011001010001",
"011000100010",
"010111110011",
"010111000101",
"010110010111",
"010101101001",
"010100111100",
"010100001111",
"010011100011",
"010010110111",
"010010001100",
"010001100001",
"010000110110",
"010000001101",
"001111100100",
"001110111011",
"001110010011",
"001101101100",
"001101000110",
"001100100000",
"001011111011",
"001011010111",
"001010110100",
"001010010001",
"001001110000",
"001001001111",
"001000101111",
"001000010000",
"000111110010",
"000111010100",
"000110111000",
"000110011101",
"000110000010",
"000101101001",
"000101010001",
"000100111010",
"000100100011",
"000100001110",
"000011111010",
"000011100111",
"000011010101",
"000011000100",
"000010110101",
"000010100110",
"000010011001",
"000010001100",
"000010000001",
"000001110111",
"000001101110",
"000001100111",
"000001100000",
"000001011011",
"000001010111",
"000001010100",
"000001010010",
"000001010001",
"000001010010",
"000001010100",
"000001010111",
"000001011011",
"000001100000",
"000001100111",
"000001101110",
"000001110111",
"000010000001",
"000010001100",
"000010011001",
"000010100110",
"000010110101",
"000011000100",
"000011010101",
"000011100111",
"000011111010",
"000100001110",
"000100100011",
"000100111010",
"000101010001",
"000101101001",
"000110000010",
"000110011101",
"000110111000",
"000111010100",
"000111110010",
"001000010000",
"001000101111",
"001001001111",
"001001110000",
"001010010001",
"001010110100",
"001011010111",
"001011111011",
"001100100000",
"001101000110",
"001101101100",
"001110010011",
"001110111011",
"001111100100",
"010000001101",
"010000110110",
"010001100001",
"010010001100",
"010010110111",
"010011100011",
"010100001111",
"010100111100",
"010101101001",
"010110010111",
"010111000101",
"010111110011",
"011000100010",
"011001010001",
"011010000000",
"011010101111",
"011011011111",
"011100001111",
"011100111111",
"011101101111",
"011110011111",
"011111001111",
"011111111111",
"100000110000",
"100001100000",
"100010010000",
"100011000000",
"100011110000",
"100100100000",
"100101010000",
"100101111111",
"100110101110",
"100111011101",
"101000001100",
"101000111010",
"101001101000",
"101010010110",
"101011000011",
"101011110000",
"101100011100",
"101101001000",
"101101110011",
"101110011110",
"101111001001",
"101111110010",
"110000011011",
"110001000100",
"110001101100",
"110010010011",
"110010111001",
"110011011111",
"110100000100",
"110100101000",
"110101001011",
"110101101110",
"110110001111",
"110110110000",
"110111010000",
"110111101111",
"111000001101",
"111000101011",
"111001000111",
"111001100010",
"111001111101",
"111010010110",
"111010101110",
"111011000101",
"111011011100",
"111011110001",
"111100000101",
"111100011000",
"111100101010",
"111100111011",
"111101001010",
"111101011001",
"111101100110",
"111101110011",
"111101111110",
"111110001000",
"111110010001",
"111110011000",
"111110011111",
"111110100100",
"111110101000",
"111110101011",
"111110101101",
"111110101110",
"111110101101",
"111110101011",
"111110101000",
"111110100100",
"111110011111",
"111110011000",
"111110010001",
"111110001000",
"111101111110",
"111101110011",
"111101100110",
"111101011001",
"111101001010",
"111100111011",
"111100101010",
"111100011000",
"111100000101",
"111011110001",
"111011011100",
"111011000101",
"111010101110",
"111010010110",
"111001111101",
"111001100010",
"111001000111",
"111000101011",
"111000001101",
"110111101111",
"110111010000",
"110110110000",
"110110001111",
"110101101110",
"110101001011",
"110100101000",
"110100000100",
"110011011111",
"110010111001",
"110010010011",
"110001101100",
"110001000100",
"110000011011",
"101111110010",
"101111001001",
"101110011110",
"101101110011",
"101101001000",
"101100011100",
"101011110000",
"101011000011",
"101010010110",
"101001101000",
"101000111010",
"101000001100",
"100111011101",
"100110101110",
"100101111111",
"100101010000",
"100100100000",
"100011110000",
"100011000000",
"100010010000",
"100001100000",
"100000110000",
"100000000000",
"011111001111",
"011110011111",
"011101101111",
"011100111111",
"011100001111",
"011011011111",
"011010101111",
"011010000000",
"011001010001",
"011000100010",
"010111110011",
"010111000101",
"010110010111",
"010101101001",
"010100111100",
"010100001111",
"010011100011",
"010010110111",
"010010001100",
"010001100001",
"010000110110",
"010000001101",
"001111100100",
"001110111011",
"001110010011",
"001101101100",
"001101000110",
"001100100000",
"001011111011",
"001011010111",
"001010110100",
"001010010001",
"001001110000",
"001001001111",
"001000101111",
"001000010000",
"000111110010",
"000111010100",
"000110111000",
"000110011101",
"000110000010",
"000101101001",
"000101010001",
"000100111010",
"000100100011",
"000100001110",
"000011111010",
"000011100111",
"000011010101",
"000011000100",
"000010110101",
"000010100110",
"000010011001",
"000010001100",
"000010000001",
"000001110111",
"000001101110",
"000001100111",
"000001100000",
"000001011011",
"000001010111",
"000001010100",
"000001010010",
"000001010001",
"000001010010",
"000001010100",
"000001010111",
"000001011011",
"000001100000",
"000001100111",
"000001101110",
"000001110111",
"000010000001",
"000010001100",
"000010011001",
"000010100110",
"000010110101",
"000011000100",
"000011010101",
"000011100111",
"000011111010",
"000100001110",
"000100100011",
"000100111010",
"000101010001",
"000101101001",
"000110000010",
"000110011101",
"000110111000",
"000111010100",
"000111110010",
"001000010000",
"001000101111",
"001001001111",
"001001110000",
"001010010001",
"001010110100",
"001011010111",
"001011111011",
"001100100000",
"001101000110",
"001101101100",
"001110010011",
"001110111011",
"001111100100",
"010000001101",
"010000110110",
"010001100001",
"010010001100",
"010010110111",
"010011100011",
"010100001111",
"010100111100",
"010101101001",
"010110010111",
"010111000101",
"010111110011",
"011000100010",
"011001010001",
"011010000000",
"011010101111",
"011011011111",
"011100001111",
"011100111111",
"011101101111",
"011110011111",
"011111001111",
"011111111111",
"100000110000",
"100001100000",
"100010010000",
"100011000000",
"100011110000",
"100100100000",
"100101010000",
"100101111111",
"100110101110",
"100111011101",
"101000001100",
"101000111010",
"101001101000",
"101010010110",
"101011000011",
"101011110000",
"101100011100",
"101101001000",
"101101110011",
"101110011110",
"101111001001",
"101111110010",
"110000011011",
"110001000100",
"110001101100",
"110010010011",
"110010111001",
"110011011111",
"110100000100",
"110100101000",
"110101001011",
"110101101110",
"110110001111",
"110110110000",
"110111010000",
"110111101111",
"111000001101",
"111000101011",
"111001000111",
"111001100010",
"111001111101",
"111010010110",
"111010101110",
"111011000101",
"111011011100",
"111011110001",
"111100000101",
"111100011000",
"111100101010",
"111100111011",
"111101001010",
"111101011001",
"111101100110",
"111101110011",
"111101111110",
"111110001000",
"111110010001",
"111110011000",
"111110011111",
"111110100100",
"111110101000",
"111110101011",
"111110101101",
"111110101110",
"111110101101",
"111110101011",
"111110101000",
"111110100100",
"111110011111",
"111110011000",
"111110010001",
"111110001000",
"111101111110",
"111101110011",
"111101100110",
"111101011001",
"111101001010",
"111100111011",
"111100101010",
"111100011000",
"111100000101",
"111011110001",
"111011011100",
"111011000101",
"111010101110",
"111010010110",
"111001111101",
"111001100010",
"111001000111",
"111000101011",
"111000001101",
"110111101111",
"110111010000",
"110110110000",
"110110001111",
"110101101110",
"110101001011",
"110100101000",
"110100000100",
"110011011111",
"110010111001",
"110010010011",
"110001101100",
"110001000100",
"110000011011",
"101111110010",
"101111001001",
"101110011110",
"101101110011",
"101101001000",
"101100011100",
"101011110000",
"101011000011",
"101010010110",
"101001101000",
"101000111010",
"101000001100",
"100111011101",
"100110101110",
"100101111111",
"100101010000",
"100100100000",
"100011110000",
"100011000000",
"100010010000",
"100001100000",
"100000110000",
"100000000000",
"011111001111",
"011110011111",
"011101101111",
"011100111111",
"011100001111",
"011011011111",
"011010101111",
"011010000000",
"011001010001",
"011000100010",
"010111110011",
"010111000101",
"010110010111",
"010101101001",
"010100111100",
"010100001111",
"010011100011",
"010010110111",
"010010001100",
"010001100001",
"010000110110",
"010000001101",
"001111100100",
"001110111011",
"001110010011",
"001101101100",
"001101000110",
"001100100000",
"001011111011",
"001011010111",
"001010110100",
"001010010001",
"001001110000",
"001001001111",
"001000101111",
"001000010000",
"000111110010",
"000111010100",
"000110111000",
"000110011101",
"000110000010",
"000101101001",
"000101010001",
"000100111010",
"000100100011",
"000100001110",
"000011111010",
"000011100111",
"000011010101",
"000011000100",
"000010110101",
"000010100110",
"000010011001",
"000010001100",
"000010000001",
"000001110111",
"000001101110",
"000001100111",
"000001100000",
"000001011011",
"000001010111",
"000001010100",
"000001010010",
"000001010001",
"000001010010",
"000001010100",
"000001010111",
"000001011011",
"000001100000",
"000001100111",
"000001101110",
"000001110111",
"000010000001",
"000010001100",
"000010011001",
"000010100110",
"000010110101",
"000011000100",
"000011010101",
"000011100111",
"000011111010",
"000100001110",
"000100100011",
"000100111010",
"000101010001",
"000101101001",
"000110000010",
"000110011101",
"000110111000",
"000111010100",
"000111110010",
"001000010000",
"001000101111",
"001001001111",
"001001110000",
"001010010001",
"001010110100",
"001011010111",
"001011111011",
"001100100000",
"001101000110",
"001101101100",
"001110010011",
"001110111011",
"001111100100",
"010000001101",
"010000110110",
"010001100001",
"010010001100",
"010010110111",
"010011100011",
"010100001111",
"010100111100",
"010101101001",
"010110010111",
"010111000101",
"010111110011",
"011000100010",
"011001010001",
"011010000000",
"011010101111",
"011011011111",
"011100001111",
"011100111111",
"011101101111",
"011110011111",
"011111001111",
"100000000000",
"100000110000",
"100001100000",
"100010010000",
"100011000000",
"100011110000",
"100100100000",
"100101010000",
"100101111111",
"100110101110",
"100111011101",
"101000001100",
"101000111010",
"101001101000",
"101010010110",
"101011000011",
"101011110000",
"101100011100",
"101101001000",
"101101110011",
"101110011110",
"101111001001",
"101111110010",
"110000011011",
"110001000100",
"110001101100",
"110010010011",
"110010111001",
"110011011111",
"110100000100",
"110100101000"
);

constant R2 : matrix_index :=(
"100000000000",
"100000110000",
"100001100000",
"100010010000",
"100011000000",
"100011110000",
"100100100000",
"100101010000",
"100101111111",
"100110101110",
"100111011101",
"101000001100",
"101000111010",
"101001101000",
"101010010110",
"101011000011",
"101011110000",
"101100011100",
"101101001000",
"101101110011",
"101110011110",
"101111001001",
"101111110010",
"110000011011",
"110001000100",
"110001101100",
"110010010011",
"110010111001",
"110011011111",
"110100000100",
"110100101000",
"110101001011",
"110101101110",
"110110001111",
"110110110000",
"110111010000",
"110111101111",
"111000001101",
"111000101011",
"111001000111",
"111001100010",
"111001111101",
"111010010110",
"111010101110",
"111011000101",
"111011011100",
"111011110001",
"111100000101",
"111100011000",
"111100101010",
"111100111011",
"111101001010",
"111101011001",
"111101100110",
"111101110011",
"111101111110",
"111110001000",
"111110010001",
"111110011000",
"111110011111",
"111110100100",
"111110101000",
"111110101011",
"111110101101",
"111110101110",
"111110101101",
"111110101011",
"111110101000",
"111110100100",
"111110011111",
"111110011000",
"111110010001",
"111110001000",
"111101111110",
"111101110011",
"111101100110",
"111101011001",
"111101001010",
"111100111011",
"111100101010",
"111100011000",
"111100000101",
"111011110001",
"111011011100",
"111011000101",
"111010101110",
"111010010110",
"111001111101",
"111001100010",
"111001000111",
"111000101011",
"111000001101",
"110111101111",
"110111010000",
"110110110000",
"110110001111",
"110101101110",
"110101001011",
"110100101000",
"110100000100",
"110011011111",
"110010111001",
"110010010011",
"110001101100",
"110001000100",
"110000011011",
"101111110010",
"101111001001",
"101110011110",
"101101110011",
"101101001000",
"101100011100",
"101011110000",
"101011000011",
"101010010110",
"101001101000",
"101000111010",
"101000001100",
"100111011101",
"100110101110",
"100101111111",
"100101010000",
"100100100000",
"100011110000",
"100011000000",
"100010010000",
"100001100000",
"100000110000",
"100000000000",
"011111001111",
"011110011111",
"011101101111",
"011100111111",
"011100001111",
"011011011111",
"011010101111",
"011010000000",
"011001010001",
"011000100010",
"010111110011",
"010111000101",
"010110010111",
"010101101001",
"010100111100",
"010100001111",
"010011100011",
"010010110111",
"010010001100",
"010001100001",
"010000110110",
"010000001101",
"001111100100",
"001110111011",
"001110010011",
"001101101100",
"001101000110",
"001100100000",
"001011111011",
"001011010111",
"001010110100",
"001010010001",
"001001110000",
"001001001111",
"001000101111",
"001000010000",
"000111110010",
"000111010100",
"000110111000",
"000110011101",
"000110000010",
"000101101001",
"000101010001",
"000100111010",
"000100100011",
"000100001110",
"000011111010",
"000011100111",
"000011010101",
"000011000100",
"000010110101",
"000010100110",
"000010011001",
"000010001100",
"000010000001",
"000001110111",
"000001101110",
"000001100111",
"000001100000",
"000001011011",
"000001010111",
"000001010100",
"000001010010",
"000001010001",
"000001010010",
"000001010100",
"000001010111",
"000001011011",
"000001100000",
"000001100111",
"000001101110",
"000001110111",
"000010000001",
"000010001100",
"000010011001",
"000010100110",
"000010110101",
"000011000100",
"000011010101",
"000011100111",
"000011111010",
"000100001110",
"000100100011",
"000100111010",
"000101010001",
"000101101001",
"000110000010",
"000110011101",
"000110111000",
"000111010100",
"000111110010",
"001000010000",
"001000101111",
"001001001111",
"001001110000",
"001010010001",
"001010110100",
"001011010111",
"001011111011",
"001100100000",
"001101000110",
"001101101100",
"001110010011",
"001110111011",
"001111100100",
"010000001101",
"010000110110",
"010001100001",
"010010001100",
"010010110111",
"010011100011",
"010100001111",
"010100111100",
"010101101001",
"010110010111",
"010111000101",
"010111110011",
"011000100010",
"011001010001",
"011010000000",
"011010101111",
"011011011111",
"011100001111",
"011100111111",
"011101101111",
"011110011111",
"011111001111",
"011111111111",
"100000110000",
"100001100000",
"100010010000",
"100011000000",
"100011110000",
"100100100000",
"100101010000",
"100101111111",
"100110101110",
"100111011101",
"101000001100",
"101000111010",
"101001101000",
"101010010110",
"101011000011",
"101011110000",
"101100011100",
"101101001000",
"101101110011",
"101110011110",
"101111001001",
"101111110010",
"110000011011",
"110001000100",
"110001101100",
"110010010011",
"110010111001",
"110011011111",
"110100000100",
"110100101000",
"110101001011",
"110101101110",
"110110001111",
"110110110000",
"110111010000",
"110111101111",
"111000001101",
"111000101011",
"111001000111",
"111001100010",
"111001111101",
"111010010110",
"111010101110",
"111011000101",
"111011011100",
"111011110001",
"111100000101",
"111100011000",
"111100101010",
"111100111011",
"111101001010",
"111101011001",
"111101100110",
"111101110011",
"111101111110",
"111110001000",
"111110010001",
"111110011000",
"111110011111",
"111110100100",
"111110101000",
"111110101011",
"111110101101",
"111110101110",
"111110101101",
"111110101011",
"111110101000",
"111110100100",
"111110011111",
"111110011000",
"111110010001",
"111110001000",
"111101111110",
"111101110011",
"111101100110",
"111101011001",
"111101001010",
"111100111011",
"111100101010",
"111100011000",
"111100000101",
"111011110001",
"111011011100",
"111011000101",
"111010101110",
"111010010110",
"111001111101",
"111001100010",
"111001000111",
"111000101011",
"111000001101",
"110111101111",
"110111010000",
"110110110000",
"110110001111",
"110101101110",
"110101001011",
"110100101000",
"110100000100",
"110011011111",
"110010111001",
"110010010011",
"110001101100",
"110001000100",
"110000011011",
"101111110010",
"101111001001",
"101110011110",
"101101110011",
"101101001000",
"101100011100",
"101011110000",
"101011000011",
"101010010110",
"101001101000",
"101000111010",
"101000001100",
"100111011101",
"100110101110",
"100101111111",
"100101010000",
"100100100000",
"100011110000",
"100011000000",
"100010010000",
"100001100000",
"100000110000",
"100000000000",
"011111001111",
"011110011111",
"011101101111",
"011100111111",
"011100001111",
"011011011111",
"011010101111",
"011010000000",
"011001010001",
"011000100010",
"010111110011",
"010111000101",
"010110010111",
"010101101001",
"010100111100",
"010100001111",
"010011100011",
"010010110111",
"010010001100",
"010001100001",
"010000110110",
"010000001101",
"001111100100",
"001110111011",
"001110010011",
"001101101100",
"001101000110",
"001100100000",
"001011111011",
"001011010111",
"001010110100",
"001010010001",
"001001110000",
"001001001111",
"001000101111",
"001000010000",
"000111110010",
"000111010100",
"000110111000",
"000110011101",
"000110000010",
"000101101001",
"000101010001",
"000100111010",
"000100100011",
"000100001110",
"000011111010",
"000011100111",
"000011010101",
"000011000100",
"000010110101",
"000010100110",
"000010011001",
"000010001100",
"000010000001",
"000001110111",
"000001101110",
"000001100111",
"000001100000",
"000001011011",
"000001010111",
"000001010100",
"000001010010",
"000001010001",
"000001010010",
"000001010100",
"000001010111",
"000001011011",
"000001100000",
"000001100111",
"000001101110",
"000001110111",
"000010000001",
"000010001100",
"000010011001",
"000010100110",
"000010110101",
"000011000100",
"000011010101",
"000011100111",
"000011111010",
"000100001110",
"000100100011",
"000100111010",
"000101010001",
"000101101001",
"000110000010",
"000110011101",
"000110111000",
"000111010100",
"000111110010",
"001000010000",
"001000101111",
"001001001111",
"001001110000",
"001010010001",
"001010110100",
"001011010111",
"001011111011",
"001100100000",
"001101000110",
"001101101100",
"001110010011",
"001110111011",
"001111100100",
"010000001101",
"010000110110",
"010001100001",
"010010001100",
"010010110111",
"010011100011",
"010100001111",
"010100111100",
"010101101001",
"010110010111",
"010111000101",
"010111110011",
"011000100010",
"011001010001",
"011010000000",
"011010101111",
"011011011111",
"011100001111",
"011100111111",
"011101101111",
"011110011111",
"011111001111",
"011111111111",
"100000110000",
"100001100000",
"100010010000",
"100011000000",
"100011110000",
"100100100000",
"100101010000",
"100101111111",
"100110101110",
"100111011101",
"101000001100",
"101000111010",
"101001101000",
"101010010110",
"101011000011",
"101011110000",
"101100011100",
"101101001000",
"101101110011",
"101110011110",
"101111001001",
"101111110010",
"110000011011",
"110001000100",
"110001101100",
"110010010011",
"110010111001",
"110011011111",
"110100000100",
"110100101000",
"110101001011",
"110101101110",
"110110001111",
"110110110000",
"110111010000",
"110111101111",
"111000001101",
"111000101011",
"111001000111",
"111001100010",
"111001111101",
"111010010110",
"111010101110",
"111011000101",
"111011011100",
"111011110001",
"111100000101",
"111100011000",
"111100101010",
"111100111011",
"111101001010",
"111101011001",
"111101100110",
"111101110011",
"111101111110",
"111110001000",
"111110010001",
"111110011000",
"111110011111",
"111110100100",
"111110101000",
"111110101011",
"111110101101",
"111110101110",
"111110101101",
"111110101011",
"111110101000",
"111110100100",
"111110011111",
"111110011000",
"111110010001",
"111110001000",
"111101111110",
"111101110011",
"111101100110",
"111101011001",
"111101001010",
"111100111011",
"111100101010",
"111100011000",
"111100000101",
"111011110001",
"111011011100",
"111011000101",
"111010101110",
"111010010110",
"111001111101",
"111001100010",
"111001000111",
"111000101011",
"111000001101",
"110111101111",
"110111010000",
"110110110000",
"110110001111",
"110101101110",
"110101001011",
"110100101000",
"110100000100",
"110011011111",
"110010111001",
"110010010011",
"110001101100",
"110001000100",
"110000011011",
"101111110010",
"101111001001",
"101110011110",
"101101110011",
"101101001000",
"101100011100",
"101011110000",
"101011000011",
"101010010110",
"101001101000",
"101000111010",
"101000001100",
"100111011101",
"100110101110",
"100101111111",
"100101010000",
"100100100000",
"100011110000",
"100011000000",
"100010010000",
"100001100000",
"100000110000",
"100000000000",
"011111001111",
"011110011111",
"011101101111",
"011100111111",
"011100001111",
"011011011111",
"011010101111",
"011010000000",
"011001010001",
"011000100010",
"010111110011",
"010111000101",
"010110010111",
"010101101001",
"010100111100",
"010100001111",
"010011100011",
"010010110111",
"010010001100",
"010001100001",
"010000110110",
"010000001101",
"001111100100",
"001110111011",
"001110010011",
"001101101100",
"001101000110",
"001100100000",
"001011111011",
"001011010111",
"001010110100",
"001010010001",
"001001110000",
"001001001111",
"001000101111",
"001000010000",
"000111110010",
"000111010100",
"000110111000",
"000110011101",
"000110000010",
"000101101001",
"000101010001",
"000100111010",
"000100100011",
"000100001110",
"000011111010",
"000011100111",
"000011010101",
"000011000100",
"000010110101",
"000010100110",
"000010011001",
"000010001100",
"000010000001",
"000001110111",
"000001101110",
"000001100111",
"000001100000",
"000001011011",
"000001010111",
"000001010100",
"000001010010",
"000001010001",
"000001010010",
"000001010100",
"000001010111",
"000001011011",
"000001100000",
"000001100111",
"000001101110",
"000001110111",
"000010000001",
"000010001100",
"000010011001",
"000010100110",
"000010110101",
"000011000100",
"000011010101",
"000011100111",
"000011111010",
"000100001110",
"000100100011",
"000100111010",
"000101010001",
"000101101001",
"000110000010",
"000110011101",
"000110111000",
"000111010100",
"000111110010",
"001000010000",
"001000101111",
"001001001111",
"001001110000",
"001010010001",
"001010110100",
"001011010111",
"001011111011",
"001100100000",
"001101000110",
"001101101100",
"001110010011",
"001110111011",
"001111100100",
"010000001101",
"010000110110",
"010001100001",
"010010001100",
"010010110111",
"010011100011",
"010100001111",
"010100111100",
"010101101001",
"010110010111",
"010111000101",
"010111110011",
"011000100010",
"011001010001",
"011010000000",
"011010101111",
"011011011111",
"011100001111",
"011100111111",
"011101101111",
"011110011111",
"011111001111",
"011111111111",
"100000110000",
"100001100000",
"100010010000",
"100011000000",
"100011110000",
"100100100000",
"100101010000",
"100101111111",
"100110101110",
"100111011101",
"101000001100",
"101000111010",
"101001101000",
"101010010110",
"101011000011",
"101011110000",
"101100011100",
"101101001000",
"101101110011",
"101110011110",
"101111001001",
"101111110010",
"110000011011",
"110001000100",
"110001101100",
"110010010011",
"110010111001",
"110011011111",
"110100000100",
"110100101000",
"110101001011",
"110101101110",
"110110001111",
"110110110000",
"110111010000",
"110111101111",
"111000001101",
"111000101011",
"111001000111",
"111001100010",
"111001111101",
"111010010110",
"111010101110",
"111011000101",
"111011011100",
"111011110001",
"111100000101",
"111100011000",
"111100101010",
"111100111011",
"111101001010",
"111101011001",
"111101100110",
"111101110011",
"111101111110",
"111110001000",
"111110010001",
"111110011000",
"111110011111",
"111110100100",
"111110101000",
"111110101011",
"111110101101",
"111110101110",
"111110101101",
"111110101011",
"111110101000",
"111110100100",
"111110011111",
"111110011000",
"111110010001",
"111110001000",
"111101111110",
"111101110011",
"111101100110",
"111101011001",
"111101001010",
"111100111011",
"111100101010",
"111100011000",
"111100000101",
"111011110001",
"111011011100",
"111011000101",
"111010101110",
"111010010110",
"111001111101",
"111001100010",
"111001000111",
"111000101011",
"111000001101",
"110111101111",
"110111010000",
"110110110000",
"110110001111",
"110101101110",
"110101001011",
"110100101000",
"110100000100",
"110011011111",
"110010111001",
"110010010011",
"110001101100",
"110001000100",
"110000011011",
"101111110010",
"101111001001",
"101110011110",
"101101110011",
"101101001000",
"101100011100",
"101011110000",
"101011000011",
"101010010110",
"101001101000",
"101000111010",
"101000001100",
"100111011101",
"100110101110",
"100101111111",
"100101010000",
"100100100000",
"100011110000",
"100011000000",
"100010010000",
"100001100000",
"100000110000",
"100000000000",
"011111001111",
"011110011111",
"011101101111",
"011100111111",
"011100001111",
"011011011111",
"011010101111",
"011010000000",
"011001010001",
"011000100010",
"010111110011",
"010111000101",
"010110010111",
"010101101001",
"010100111100",
"010100001111",
"010011100011",
"010010110111",
"010010001100",
"010001100001",
"010000110110",
"010000001101",
"001111100100",
"001110111011",
"001110010011",
"001101101100",
"001101000110",
"001100100000",
"001011111011",
"001011010111",
"001010110100",
"001010010001",
"001001110000",
"001001001111",
"001000101111",
"001000010000",
"000111110010",
"000111010100",
"000110111000",
"000110011101",
"000110000010",
"000101101001",
"000101010001",
"000100111010",
"000100100011",
"000100001110",
"000011111010",
"000011100111",
"000011010101",
"000011000100",
"000010110101",
"000010100110",
"000010011001",
"000010001100",
"000010000001",
"000001110111",
"000001101110",
"000001100111",
"000001100000",
"000001011011",
"000001010111",
"000001010100",
"000001010010",
"000001010001",
"000001010010",
"000001010100",
"000001010111",
"000001011011",
"000001100000",
"000001100111",
"000001101110",
"000001110111",
"000010000001",
"000010001100",
"000010011001",
"000010100110",
"000010110101",
"000011000100",
"000011010101",
"000011100111",
"000011111010",
"000100001110",
"000100100011",
"000100111010",
"000101010001",
"000101101001",
"000110000010",
"000110011101",
"000110111000",
"000111010100",
"000111110010",
"001000010000",
"001000101111",
"001001001111",
"001001110000",
"001010010001",
"001010110100",
"001011010111",
"001011111011",
"001100100000",
"001101000110",
"001101101100",
"001110010011",
"001110111011",
"001111100100",
"010000001101",
"010000110110",
"010001100001",
"010010001100",
"010010110111",
"010011100011",
"010100001111",
"010100111100",
"010101101001",
"010110010111",
"010111000101",
"010111110011",
"011000100010",
"011001010001",
"011010000000",
"011010101111",
"011011011111",
"011100001111",
"011100111111",
"011101101111",
"011110011111",
"011111001111"
);

begin
number <= conv_integer (num);
process(clk)
begin
if (CLK'EVENT and CLK = '1') then
    da1 <= R1(number);
    da2 <= R2(number);
end if;
end process;

end Behavioral;

